library verilog;
use verilog.vl_types.all;
entity ej_a_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ej_a_vlg_check_tst;
