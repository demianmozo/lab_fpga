library verilog;
use verilog.vl_types.all;
entity ej_a_vlg_vec_tst is
end ej_a_vlg_vec_tst;
